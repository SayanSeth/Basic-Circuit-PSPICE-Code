Common Base Amplifier
Vs 6 0 AC 1 SIN(0 10M 1KHZ)
VCC 5 0 DC 12
R1 5 4 1.2K
R2 5 3 22K
R3 2 0 220
R4 3 0 3.3K
C1 3 0 1U
C2 4 7 1U
C3 2 6 1U
RL 7 0 100K
Q1 4 3 2 BC107b

.model BC107b   NPN (IS =1.8E-14 ISE=5.0E-14 NF =.9955 NE =1.46
+					 BF =200 BR =35.5 IKF=.14 IKR=.03 ISC=1.72E-13
+					 NC =1.27 NR =1.005 RB =.56 RE =.6 RC =.25 VAF=80
+					 VAR=12.5 CJE=13E-12 TF =.64E-9 CJC=4E-12 TR =50.72E-9
+					 VJC=.54 MJC=.33)
*
* ANALYSIS
.AC DEC 5 10 1000MEG
*.OP
*.TRAN 0 5M
.END
