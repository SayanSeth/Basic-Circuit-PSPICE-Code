RC Coupled Amplifier
VS 8 0 AC 1 SIN(0 10M 1KHZ)
VCC 1 0 DC 12
R1 1 4 1k
R2 1 2 1k
R3 3 0 1k
R4 2 0 1k
R5 7 0 1k
R6 5 0 1k
R7 6 1 1k
R8 5 1 1k
C1 3 0 1u
C2 7 0 1u
C3 4 5 1u
C4 8 2 1u
C5 6 9 1u
RL 9 0 100k
Q2 6 5 7 BC107b
Q1 4 2 3 BC107b

.model BC107b   NPN(IS =1.8E-14 ISE=5.0E-14 NF =.9955 NE =1.46
+				BF =200 BR =35.5 IKF=.14 IKR=.03 ISC=1.72E-13 NC =1.27 NR =1.005
+				RB =.56 RE =.6 RC =.25 VAF=80 VAR=12.5 CJE=13E-12 TF =.64E-9 CJC=4E-12
+				TR =50.72E-9 VJC=.54 MJC=.33)
*
* ANALYSIS
*.AC DEC 5 1 1000MEG
*.OP
*.PROBE
.TRAN 0.5M 5M
.END
